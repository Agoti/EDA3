library verilog;
use verilog.vl_types.all;
entity Buzzer_vlg_vec_tst is
end Buzzer_vlg_vec_tst;
